module main;
  initial 
    begin
      $display("2022");
      $display("01");
      $display("08");
      $finish ;
    end
endmodule
